module drive_dac
(
	input  [9:0] sw,
	output [40:0] gpio1,
	output  [9:0] led
); 

	//assign led = sw;
	
endmodule