library verilog;
use verilog.vl_types.all;
entity deserializer_vlg_vec_tst is
end deserializer_vlg_vec_tst;
